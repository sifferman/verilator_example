module test;
    initial $display("Hello");
endmodule
